////
//
// University of Utah ECE 5710/6710 Edge Detection ASIC
//
// Create Date: 10/23/2020
// Module Name: colorspace_converter
// Description: Converts an RGB colorspace input to grayscale.
// Authors: Jacob Peterson
//
////

module colorspace_converter();

endmodule

////
//
// University of Utah ECE 5710/6710 Edge Detection ASIC
//
// Create Date: 10/28/2020
// Module Name: buffered_matrix_colorspace_converter
// Description: Converts an RGB colorspace VGA input to a grayscaled pixel matrix output.
// Authors: Jacob Peterson
//
////

module buffered_matrix3_colorspace_converter
    #(
    parameter integer P_FRAME_COLUMNS = 640, // The number of columns in the frame
    parameter integer P_FRAME_ROWS = 480, // The number of rows in the frame
    parameter integer P_PIXEL_DEPTH = 24, // The color depth of the pixel (MUST be a multiple of 3)

    // START port list local parameters

    parameter integer P_FRAME_COLUMN_BITS = $clog2(P_FRAME_COLUMNS),
    parameter integer P_FRAME_ROW_BITS = $clog2(P_FRAME_ROWS),
    parameter integer P_SUBPIXEL_DEPTH = P_PIXEL_DEPTH / 3,

    // This is the dimension size of the square 2D pixel matrix output.
    parameter integer P_OUTPUT_MATRIX_SIZE = 3,

    // The output matrix excludes the center grayscaled pixel so we subtract one P_SUBPIXEL_DEPTH.
    parameter integer P_PIXEL_MATRIX_BITS = (P_SUBPIXEL_DEPTH * P_OUTPUT_MATRIX_SIZE * P_OUTPUT_MATRIX_SIZE) - P_SUBPIXEL_DEPTH

    // END port list local parameters
    )
    (
    input wire I_CLK, // Clock input
    input wire I_RESET, // Reset input

    input wire I_PIXEL_CLK, // Pixel clock input
    input wire I_DATA_VALID, // The data valid input (should be asserted when in the active region of the frame)
    input wire I_VSYNC, // The Vertical Sync input
    input wire [P_PIXEL_DEPTH - 1 : 0] I_PIXEL,  // RGB pixel input

    output wire [P_FRAME_COLUMN_BITS - 1 : 0] O_PIXEL_COLUMN, // The start column of the output matrix relative to the start column of the frame output
    output wire [P_FRAME_ROW_BITS - 1 : 0] O_PIXEL_ROW, // The start row of the output matrix relative to the start row of the frame output

    // The grayscaled pixel matrix output (excludes the center pixel for Sobel filter specification)
    // Format:
    // {top_left,    top,    top_right,
    //  middle_left, 	      middle_right,
    //  bottom_left, bottom, bottom_right}
    output wire [P_PIXEL_MATRIX_BITS - 1 : 0] O_PIXEL_MATRIX,
    output wire O_PIXEL_MATRIX_READY // Matrix ready output (asserted if outputs are ready/valid)
    );

    // START local parameters
    localparam P_FRAME_BUFFER_ROWS = 3; // The number of rows to use for the internal grayscaled pixel buffer
    localparam P_FRAME_BUFFER_REQUIRED_ROWS = 2; // The minimum number of rows required for a valid pixel matrix output
    localparam P_FRAME_BUFFER_REQUIRED_COLUMNS = 3; // The minimum number of columns required for a valid pixel matrix output
    // END local parameters

    // START registers and wires

    // States for input frame (synchronized with pixel clock)
    reg q_frame_column_reset; // The current state of if current frame column should be reset to zero
    wire n_frame_column_reset; // The next state of if current frame column should be reset to zero
    reg q_frame_row_reset; // The current state of if current frame row should be reset to zero
    wire n_frame_row_reset; // The next state of if current frame row should be reset to zero
    reg q_frame_row_increment_pulse; // The current state of the assertion pulse if current frame row should be incremented
    wire n_frame_row_increment_pulse; // The next state of the assertion pulse if current frame row should be incremented
    reg [P_FRAME_COLUMN_BITS - 1 : 0] q_frame_column; // The current state of the current frame pixel column
    wire [P_FRAME_COLUMN_BITS - 1 : 0] n_frame_column; // The next state of the current frame pixel column
    reg [P_FRAME_ROW_BITS - 1 : 0] q_frame_row; // The current state of the current frame pixel row
    wire [P_FRAME_ROW_BITS - 1 : 0] n_frame_row; // The next state of the current frame pixel row

    // States for iGrayscale
    wire [P_SUBPIXEL_DEPTH - 1 : 0] grayscaled_pixel; // Grayscale output of the directly-inputted pixel

    // States for iGrayscaledFrameBufferMatrix3
    wire should_frame_buffer_increment; // Asserted if the frame buffer should start counting in sync with the input pixel clock
    reg q_frame_buffer_column_reset; // The current state of if current frame buffer column should be reset to zero
    wire n_frame_buffer_column_reset; // The next state of if current frame buffer column should be reset to zero
    reg q_frame_buffer_row_reset; // The current state of if current frame buffer row should be reset to zero
    wire n_frame_buffer_row_reset; // The next state of if current frame buffer row should be reset to zero
    reg q_frame_buffer_row_increment_pulse; // The current state of the assertion pulse if current frame buffer row should be incremented
    wire n_frame_buffer_row_increment_pulse; // The next state of the assertion pulse if current frame buffer row should be incremented
    reg [P_FRAME_COLUMN_BITS - 1 : 0] q_frame_buffer_column; // The current state of the frame buffer column index
    wire [P_FRAME_COLUMN_BITS - 1 : 0] n_frame_buffer_column; // The next state of the frame buffer column index
    reg [P_FRAME_ROW_BITS - 1 : 0] q_frame_buffer_row; // The current state of the frame buffer row index
    wire [P_FRAME_ROW_BITS - 1 : 0] n_frame_buffer_row; // The next state of the frame buffer row index
    reg q_frame_buffer_write_enable; // The current state of if the frame buffer should enable writing
    wire n_frame_buffer_write_enable; // The next state of if the frame buffer should enable writing
    reg q_frame_buffer_read_enable; // The current state of if the frame buffer should enable reading
    wire n_frame_buffer_read_enable; // The next state of if the frame buffer should enable reading

    // States for logic
    reg q_frame_buffer_write_pulse; // The current state of the assertion pulse if the buffered should be written to
    wire n_frame_buffer_write_pulse; // The next state of the assertion pulse if the buffered should be written to

    // States for output
    reg [P_FRAME_COLUMN_BITS - 1 : 0] q_o_pixel_column; // The current state of the output pixel column
    wire [P_FRAME_COLUMN_BITS - 1 : 0] n_o_pixel_column; // The next state of the output pixel column
    reg [P_FRAME_ROW_BITS - 1 : 0] q_o_pixel_row; // The current state of the output pixel row
    wire [P_FRAME_ROW_BITS - 1 : 0] n_o_pixel_row; // The next state of the output pixel row
    reg [P_PIXEL_MATRIX_BITS - 1 : 0] q_o_pixel_matrix; // The current state of the output pixel matrix
    wire [P_PIXEL_MATRIX_BITS - 1 : 0] n_o_pixel_matrix; // The next state of the output pixel matrix
    reg q_o_pixel_matrix_ready; // The current state of the output pixel matrix ready signal
    wire n_o_pixel_matrix_ready; // The next state of the output pixel matrix ready signal

    // END registers and wires

    // START output mapping
    assign O_PIXEL_COLUMN = q_o_pixel_column;
    assign O_PIXEL_ROW = q_o_pixel_row;
    assign O_PIXEL_MATRIX = q_o_pixel_matrix;
    assign O_PIXEL_MATRIX_READY = q_o_pixel_matrix_ready;
    // END output mapping

    // START RTL logic
    assign n_frame_column_reset = ~I_DATA_VALID;
    assign n_frame_row_reset = ~I_VSYNC;
    assign n_frame_row_increment_pulse = I_DATA_VALID ? 1'b0 : (q_frame_row_increment_pulse ? 1'b0 : 1'b1);
    assign n_frame_column = q_frame_column_reset ? {P_FRAME_COLUMN_BITS{1'b0}} : q_frame_column + 1'b1;
    assign n_frame_row = q_frame_row_reset ? {P_FRAME_ROW_BITS{1'b0}} :
                (q_frame_row_increment_pulse ? q_frame_row + 1'b1 : q_frame_row);

    assign should_frame_buffer_increment = q_frame_column >= P_FRAME_BUFFER_REQUIRED_COLUMNS - 1 &&
                q_frame_row >= P_FRAME_BUFFER_REQUIRED_ROWS - 1;

    assign n_frame_buffer_column_reset = ~I_DATA_VALID;
    assign n_frame_buffer_row_reset = ~I_VSYNC;
    assign n_frame_buffer_row_increment_pulse = I_DATA_VALID ? 1'b0 : (q_frame_buffer_row_increment_pulse ? 1'b0 : 1'b1);
    assign n_frame_buffer_column = q_frame_buffer_column_reset ? {P_FRAME_COLUMN_BITS{1'b0}} : q_frame_buffer_column + 1'b1;
    assign n_frame_buffer_row = q_frame_buffer_row_reset ? {P_FRAME_ROW_BITS{1'b0}} :
                (q_frame_buffer_row_increment_pulse ? q_frame_buffer_row + 1'b1 : q_frame_buffer_row);
    // END RTL logic

    // START module instantiations
    grayscale #(
        .P_PIXEL_DEPTH(P_PIXEL_DEPTH)
        )
        iGrayscale
        (
        .I_CLK(I_CLK),
        .I_RESET(I_RESET),
        .I_PIXEL(I_PIXEL),

        .O_PIXEL(grayscaled_pixel)
        );

    frame_buffer_matrix3 #(
        .P_COLUMNS(P_FRAME_COLUMNS),
        .P_ROWS(P_FRAME_BUFFER_ROWS),
        .P_PIXEL_DEPTH(P_SUBPIXEL_DEPTH)
        )
        iGrayscaledFrameBufferMatrix3
        (
        .I_CLK(I_CLK),
        .I_RESET(I_RESET),
        .I_COLUMN(q_frame_buffer_column),
        .I_ROW(q_frame_buffer_row),
        .I_PIXEL(grayscaled_pixel),
        .I_WRITE_ENABLE(q_frame_buffer_write_enable),
        .I_READ_ENABLE(q_frame_buffer_read_enable),

        .O_PIXEL_MATRIX(n_o_pixel_matrix)
        );
    // END module instantiations

    // Clock block
    always @(posedge I_CLK) begin
        if (I_RESET) begin
            q_frame_buffer_column <= {P_FRAME_COLUMN_BITS{1'b0}};
            q_frame_buffer_row <= {P_FRAME_ROW_BITS{1'b0}};
            q_frame_buffer_write_enable <= 1'b0;
            q_frame_buffer_read_enable <= 1'b0;

            q_frame_buffer_write_pulse <= 1'b0;

            q_o_pixel_column <= {P_FRAME_COLUMN_BITS{1'b0}};
            q_o_pixel_row <= {P_FRAME_ROW_BITS{1'b0}};
            q_o_pixel_matrix <= {P_PIXEL_MATRIX_BITS{1'b0}};
            q_o_pixel_matrix_ready <= 1'b0;
        end else begin
            q_frame_buffer_column <= n_frame_buffer_column;
            q_frame_buffer_row <= n_frame_buffer_row;
            q_frame_buffer_write_enable <= n_frame_buffer_write_enable;
            q_frame_buffer_read_enable <= n_frame_buffer_read_enable;

            q_frame_buffer_write_pulse <= n_frame_buffer_write_pulse;

            q_o_pixel_column <= n_o_pixel_column;
            q_o_pixel_row <= n_o_pixel_row;
            q_o_pixel_matrix <= n_o_pixel_matrix;
            q_o_pixel_matrix_ready <= n_o_pixel_matrix_ready;
        end
    end

    // Pixel clock block
    always @(posedge I_PIXEL_CLK) begin
        if (I_RESET) begin
            q_frame_column_reset <= 1'b0;
            q_frame_row_reset <= 1'b0;
            q_frame_row_increment_pulse <= 1'b0;
            q_frame_column <= {P_FRAME_COLUMN_BITS{1'b0}};
            q_frame_row <= {P_FRAME_ROW_BITS{1'b0}};

            q_frame_buffer_column_reset <= 1'b0;
            q_frame_buffer_row_reset <= 1'b0;
            q_frame_buffer_row_increment_pulse <= 1'b0;
            q_frame_buffer_column <= {P_FRAME_COLUMN_BITS{1'b0}};
            q_frame_buffer_row <= {P_FRAME_ROW_BITS{1'b0}};
        end else begin
            q_frame_column_reset <= n_frame_column_reset;
            q_frame_row_reset <= n_frame_row_reset;
            q_frame_row_increment_pulse <= n_frame_row_increment_pulse;
            q_frame_column <= n_frame_column;
            q_frame_row <= n_frame_row;

            q_frame_buffer_column_reset <= n_frame_buffer_column_reset;
            q_frame_buffer_row_reset <= n_frame_buffer_row_reset;
            q_frame_buffer_row_increment_pulse <= n_frame_buffer_row_increment_pulse;
            q_frame_buffer_column <= n_frame_buffer_column;
            q_frame_buffer_row <= n_frame_buffer_row;
        end
    end
endmodule

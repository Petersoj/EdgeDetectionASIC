////
//
// University of Utah ECE 5710/6710 Edge Detection ASIC
//
// Create Date: 10/23/2020
// Module Name: frame_buffer
// Description: A memory buffer for a video frame.
// Authors: Jacob Peterson
//
////

module frame_buffer();

endmodule
